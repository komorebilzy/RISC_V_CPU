`include "defines.v"
module reg_file(
    //from rob
    input wire rs1_sgn
);
endmodule